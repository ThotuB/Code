library verilog;
use verilog.vl_types.all;
entity pat_tb is
end pat_tb;
